// Reference functions that use Bluespec's '*' operator
function Bit#(TAdd#(n, n)) multiply_unsigned(Bit#(n) a, Bit#(n) b);
    UInt#(n) a_uint = unpack(a);
    UInt#(n) b_uint = unpack(b);
    UInt#(TAdd#(n, n)) product_uint = zeroExtend(a_uint) * zeroExtend(b_uint);
    return pack(product_uint);
endfunction

function Bit#(TAdd#(n, n)) multiply_signed(Bit#(n) a, Bit#(n) b);
    Int#(n) a_int = unpack(a);
    Int#(n) b_int = unpack(b);
    Int#(TAdd#(n, n)) product_int = signExtend(a_int) * signExtend(b_int);
    return pack(product_int);
endfunction

// Exercise 2
// Multiplication by repeated addition
function Bit#(TAdd#(n, n)) multiply_by_adding(Bit#(n) a, Bit#(n) b);
    // silly version
    // Bit#(TAdd#(n, n)) out = '0;
    // Bit#(TAdd#(n, n)) extended_b = zeroExtend(b);
    // for (Bit#(n) i = 0; i < a; i = i + 1) begin
    //     out = out + extended_b;
    // end
    // return out;

    Bit#(TAdd#(n, n)) product = '0;
    for (Integer i = 0; i < valueOf(n); i = i + 1) begin
        // not best solution
        product = product + (zeroExtend(unpack(a[i]) ? b : '0) << i);
    end
    return product;
endfunction

// Multiplier Interface
interface Multiplier#(numeric type n);
    method Bool start_ready();
    method Action start(Bit#(n) a, Bit#(n) b);
    method Bool result_ready();
    method ActionValue#(Bit#(TAdd#(n, n))) result();
endinterface


// Exercise 4
// Folded multiplier by repeated addition
module mkFoldedMultiplier(Multiplier#(n));
endmodule



function Bit#(n) arth_shift(Bit#(n) a, Integer n, Bool right_shift);
    Int#(n) a_int = unpack(a);
    Bit#(n) out = 0;
    if (right_shift) begin
        out = pack(a_int >> n);
    end
    else begin //left shift
        out = pack(a_int << n); end
    return out;
endfunction



// Exercise 6
// Booth Multiplier
module mkBoothMultiplier(Multiplier#(n));
endmodule



// Exercise 8
// Radix-4 Booth Multiplier
module mkBoothMultiplierRadix4(Multiplier#(n));
endmodule
